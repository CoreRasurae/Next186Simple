//Copyright (C)2014-2023 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8.11 Education
//Part Number: GW2AR-LV18QN88C8/I7
//Device: GW2AR-18
//Device Version: C
//Created Time: Tue Jun 27 20:26:32 2023

module Gowin_DPB_VGAFont (douta, doutb, clka, ocea, cea, reseta, wrea, clkb, oceb, ceb, resetb, wreb, ada, dina, adb, dinb);

output [7:0] douta;
output [7:0] doutb;
input clka;
input ocea;
input cea;
input reseta;
input wrea;
input clkb;
input oceb;
input ceb;
input resetb;
input wreb;
input [11:0] ada;
input [7:0] dina;
input [11:0] adb;
input [7:0] dinb;

wire [11:0] dpb_inst_0_douta_w;
wire [11:0] dpb_inst_0_doutb_w;
wire [11:0] dpb_inst_1_douta_w;
wire [11:0] dpb_inst_1_doutb_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

DPB dpb_inst_0 (
    .DOA({dpb_inst_0_douta_w[11:0],douta[3:0]}),
    .DOB({dpb_inst_0_doutb_w[11:0],doutb[3:0]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,gw_gnd}),
    .BLKSELB({gw_gnd,gw_gnd,gw_gnd}),
    .ADA({ada[11:0],gw_gnd,gw_gnd}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[3:0]}),
    .ADB({adb[11:0],gw_gnd,gw_gnd}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[3:0]})
);

defparam dpb_inst_0.READ_MODE0 = 1'b0;
defparam dpb_inst_0.READ_MODE1 = 1'b0;
defparam dpb_inst_0.WRITE_MODE0 = 2'b00;
defparam dpb_inst_0.WRITE_MODE1 = 2'b00;
defparam dpb_inst_0.BIT_WIDTH_0 = 4;
defparam dpb_inst_0.BIT_WIDTH_1 = 4;
defparam dpb_inst_0.BLK_SEL_0 = 3'b000;
defparam dpb_inst_0.BLK_SEL_1 = 3'b000;
defparam dpb_inst_0.RESET_MODE = "SYNC";
defparam dpb_inst_0.INIT_RAM_00 = 256'h000008CEEEEC00000000EFF7BFFBFE000000E11951151E000000000000000000;
defparam dpb_inst_0.INIT_RAM_01 = 256'h0000008CC80000000000C88EFFEC80000000C88777CC80000000008CEC800000;
defparam dpb_inst_0.INIT_RAM_02 = 256'h00008CCCC8AE6E00FFFFF39DD93FFFFF00000C6226C00000FFFFFF7337FFFFFF;
defparam dpb_inst_0.INIT_RAM_03 = 256'h000088BC7CB8800000006773333F3F0000000000000F3F00000088E8C6666C00;
defparam dpb_inst_0.INIT_RAM_04 = 256'h0000660666666600000008CE888EC800000026EEEEEEE620000000008E800000;
defparam dpb_inst_0.INIT_RAM_05 = 256'h0000E8CE888EC8000000EEEE00000000000C6C8C66C806C00000BBBBBBBBBF00;
defparam dpb_inst_0.INIT_RAM_06 = 256'h00000000E00000000000008CEC80000000008CE88888880000008888888EC800;
defparam dpb_inst_0.INIT_RAM_07 = 256'h00000088CCEE000000000EECC88000000000008CEC800000000000E000000000;
defparam dpb_inst_0.INIT_RAM_08 = 256'h0000CCECCCECC00000000000000466600000880888CCC8000000000000000000;
defparam dpb_inst_0.INIT_RAM_09 = 256'h000000000000000000006CCCC68CC800000066008C6200000088C6666C026C88;
defparam dpb_inst_0.INIT_RAM_0A = 256'h00000088E88000000000006CFC600000000008CCCCCC80000000C80000008C00;
defparam dpb_inst_0.INIT_RAM_0B = 256'h000000008C620000000088000000000000000000E00000000000888000000000;
defparam dpb_inst_0.INIT_RAM_0C = 256'h0000C6666C666C000000E60008C66C000000E8888888880000008C666666C800;
defparam dpb_inst_0.INIT_RAM_0D = 256'h000000008C666E000000C6666C0008000000C6666C000E000000ECCCECCCCC00;
defparam dpb_inst_0.INIT_RAM_0E = 256'h0000088000880000000008800088000000008C666E666C000000C6666C666C00;
defparam dpb_inst_0.INIT_RAM_0F = 256'h0000880888C66C000000008C6C8000000000000E00E0000000006C80008C6000;
defparam dpb_inst_0.INIT_RAM_10 = 256'h0000C62000026C000000C6666C666C0000006666E66C80000000C0CEEE66C000;
defparam dpb_inst_0.INIT_RAM_11 = 256'h0000A666E0026C000000000088826E000000E62088826E0000008C666666C800;
defparam dpb_inst_0.INIT_RAM_12 = 256'h0000666C88C6660000008CCCCCCCCE000000C88888888C00000066666E666600;
defparam dpb_inst_0.INIT_RAM_13 = 256'h0000C66666666C0000006666EEE666000000666666EEE6000000E62000000000;
defparam dpb_inst_0.INIT_RAM_14 = 256'h0000C666C8066C0000006666CC666C0000ECCE6666666C00000000000C666C00;
defparam dpb_inst_0.INIT_RAM_15 = 256'h0000CEE666666600000008C6666666000000C666666666000000C888888AEE00;
defparam dpb_inst_0.INIT_RAM_16 = 256'h0000C00000000C000000E62008C66E000000C8888C666600000066CC88CC6600;
defparam dpb_inst_0.INIT_RAM_17 = 256'h00F00000000000000000000000006C800000CCCCCCCCCC00000026EC80000000;
defparam dpb_inst_0.INIT_RAM_18 = 256'h0000C60006C000000000C6666C80000000006CCCCC8000000000000000000800;
defparam dpb_inst_0.INIT_RAM_19 = 256'h08CCCCCCCC600000000000000004C8000000C600E6C0000000006CCCCCCCCC00;
defparam dpb_inst_0.INIT_RAM_1A = 256'h000066C88C6000000C66666666E066000000C888888088000000666666C00000;
defparam dpb_inst_0.INIT_RAM_1B = 256'h0000C66666C000000000666666C00000000066666EC000000000C88888888800;
defparam dpb_inst_0.INIT_RAM_1C = 256'h0000C6C806C000000000000066C000000ECCCCCCCC6000000000C66666C00000;
defparam dpb_inst_0.INIT_RAM_1D = 256'h0000CE666660000000008C666660000000006CCCCCC000000000C60000C00000;
defparam dpb_inst_0.INIT_RAM_1E = 256'h0000E88880888E000000E6008CE0000008C6E6666660000000006C888C600000;
defparam dpb_inst_0.INIT_RAM_1F = 256'h00000E666C800000000000000000C600000008888E8880000000888880888800;
defparam dpb_inst_0.INIT_RAM_20 = 256'h00006CCCCC80C8000000C600E6C008C000006CCCCCC00C0000C6CC6200026C00;
defparam dpb_inst_0.INIT_RAM_21 = 256'h000C6CC6006C000000006CCCCC808C8000006CCCCC80800000006CCCCC800C00;
defparam dpb_inst_0.INIT_RAM_22 = 256'h0000C888888006000000C600E6C080000000C600E6C006000000C600E6C0C800;
defparam dpb_inst_0.INIT_RAM_23 = 256'h0000666E66C808C80000666E66C800600000C888888080000000C88888806C80;
defparam dpb_inst_0.INIT_RAM_24 = 256'h0000C66666C0C8000000ECCCCECCCE000000E88E66C000000000E600C06E0008;
defparam dpb_inst_0.INIT_RAM_25 = 256'h00006CCCCCC0800000006CCCCCC0C8000000C66666C080000000C66666C00600;
defparam dpb_inst_0.INIT_RAM_26 = 256'h000088C60006C8800000C666666660600000C6666666C06008C6E66666600600;
defparam dpb_inst_0.INIT_RAM_27 = 256'h000888888E888BE000006CCCEC48CC800000888E8E8C66000000C60000004C80;
defparam dpb_inst_0.INIT_RAM_28 = 256'h00006CCCCCC000800000C66666C000800000C888888008C000006CCCCC800080;
defparam dpb_inst_0.INIT_RAM_29 = 256'h000000000C08CC80000000000E0ECCC00000666EEE6660C60000666666C0C600;
defparam dpb_inst_0.INIT_RAM_2A = 256'h00E8C6C008C62000000006666E000000000000000E0000000000C66000000000;
defparam dpb_inst_0.INIT_RAM_2B = 256'h0000008C6C8000000000006C8C60000000008CCC888088000066EEE608C62000;
defparam dpb_inst_0.INIT_RAM_2C = 256'h88888888888888887D7D7D7D7D7D7D7DA5A5A5A5A5A5A5A54141414141414141;
defparam dpb_inst_0.INIT_RAM_2D = 256'h66666666E0000000666666666666666688888888888888888888888888888888;
defparam dpb_inst_0.INIT_RAM_2E = 256'h6666666666E00000666666666666666666666666666666668888888888800000;
defparam dpb_inst_0.INIT_RAM_2F = 256'h8888888880000000000000008888888800000000E666666600000000E6666666;
defparam dpb_inst_0.INIT_RAM_30 = 256'h88888888F888888888888888F000000000000000F888888800000000F8888888;
defparam dpb_inst_0.INIT_RAM_31 = 256'h666666667666666688888888F8F8888888888888F888888800000000F0000000;
defparam dpb_inst_0.INIT_RAM_32 = 256'h6666666670F0000000000000F07666666666666670F0000000000000F0766666;
defparam dpb_inst_0.INIT_RAM_33 = 256'h00000000F0F88888666666667076666600000000F0F000006666666670766666;
defparam dpb_inst_0.INIT_RAM_34 = 256'h00000000F666666666666666F000000088888888F0F0000000000000F6666666;
defparam dpb_inst_0.INIT_RAM_35 = 256'h66666666F666666666666666F000000088888888F8F0000000000000F8F88888;
defparam dpb_inst_0.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFF88888888F0000000000000008888888888888888F8F88888;
defparam dpb_inst_0.INIT_RAM_37 = 256'h000000000FFFFFFFFFFFFFFFFFFFFFFF0000000000000000FFFFFFFFF0000000;
defparam dpb_inst_0.INIT_RAM_38 = 256'h0000CCCCCCCE00000000000000066E000000C666C8CCC80000006C888C600000;
defparam dpb_inst_0.INIT_RAM_39 = 256'h0000888888C60000000000C6666600000000088888E000000000E6008006E000;
defparam dpb_inst_0.INIT_RAM_3A = 256'h0000C6666EC80E000000ECCCC666C80000008C66E66C80000000E8C666C8E000;
defparam dpb_inst_0.INIT_RAM_3B = 256'h000066666666C0000000C0000C000C00000000E3BBE63000000000EBBBE00000;
defparam dpb_inst_0.INIT_RAM_3C = 256'h0000E0C80008C0000000E008C6C800000000F0088E88000000000E00E00E0000;
defparam dpb_inst_0.INIT_RAM_3D = 256'h000000C60C60000000000880E0880000000008888888888888888888888BBE00;
defparam dpb_inst_0.INIT_RAM_3E = 256'h0000CCCCCCCCCCF000000008000000000000000880000000000000000008CC80;
defparam dpb_inst_0.INIT_RAM_3F = 256'h000000000000000000000CCCCCCC00000000000008800800000000000CCCCC80;

DPB dpb_inst_1 (
    .DOA({dpb_inst_1_douta_w[11:0],douta[7:4]}),
    .DOB({dpb_inst_1_doutb_w[11:0],doutb[7:4]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,gw_gnd}),
    .BLKSELB({gw_gnd,gw_gnd,gw_gnd}),
    .ADA({ada[11:0],gw_gnd,gw_gnd}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[7:4]}),
    .ADB({adb[11:0],gw_gnd,gw_gnd}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[7:4]})
);

defparam dpb_inst_1.READ_MODE0 = 1'b0;
defparam dpb_inst_1.READ_MODE1 = 1'b0;
defparam dpb_inst_1.WRITE_MODE0 = 2'b00;
defparam dpb_inst_1.WRITE_MODE1 = 2'b00;
defparam dpb_inst_1.BIT_WIDTH_0 = 4;
defparam dpb_inst_1.BIT_WIDTH_1 = 4;
defparam dpb_inst_1.BLK_SEL_0 = 3'b000;
defparam dpb_inst_1.BLK_SEL_1 = 3'b000;
defparam dpb_inst_1.RESET_MODE = "SYNC";
defparam dpb_inst_1.INIT_RAM_00 = 256'h0000137FFFF6000000007FFEDFFDF70000007889A88A87000000000000000000;
defparam dpb_inst_1.INIT_RAM_01 = 256'h000000133100000000003117FF7310000000311EEE33100000000137F7310000;
defparam dpb_inst_1.INIT_RAM_02 = 256'h00007CCCC7100100FFFFFC9BB9CFFFFF0000036446300000FFFFFFECCEFFFFFF;
defparam dpb_inst_1.INIT_RAM_03 = 256'h000011D3E3D11000000CEE66666767000000EF73333333000000117136666300;
defparam dpb_inst_1.INIT_RAM_04 = 256'h00006606666666000000013711173100000000013F31000000008CEFFFFFEC80;
defparam dpb_inst_1.INIT_RAM_05 = 256'h00007137111731000000FFFF000000000007C036CC636C700000111117DDD700;
defparam dpb_inst_1.INIT_RAM_06 = 256'h00000036F630000000000010F010000000001371111111000000111111173100;
defparam dpb_inst_1.INIT_RAM_07 = 256'h0000013377FF000000000FF77331000000000026F6200000000000FCCC000000;
defparam dpb_inst_1.INIT_RAM_08 = 256'h000066F666F66000000000000002666000001101113331000000000000000000;
defparam dpb_inst_1.INIT_RAM_09 = 256'h000000000006333000007CCCD736630000008C6310CC000000117C8007CCC711;
defparam dpb_inst_1.INIT_RAM_0A = 256'h000000117110000000000063F360000000003100000013000000013333331000;
defparam dpb_inst_1.INIT_RAM_0B = 256'h00008C6310000000000011000000000000000000F00000000003111000000000;
defparam dpb_inst_1.INIT_RAM_0C = 256'h00007C000300C7000000FCC63100C7000000711111173100000036CCDDCC6300;
defparam dpb_inst_1.INIT_RAM_0D = 256'h000033331000CF0000007CCCCFCC630000007C000FCCCF0000001000FC631000;
defparam dpb_inst_1.INIT_RAM_0E = 256'h000031100011000000000110001100000000700007CCC70000007CCCC7CCC700;
defparam dpb_inst_1.INIT_RAM_0F = 256'h00001101110CC700000063100013600000000007007000000000001363100000;
defparam dpb_inst_1.INIT_RAM_10 = 256'h000036CCCCCC63000000F66667666F000000CCCCFCC6310000007CDDDDCC7000;
defparam dpb_inst_1.INIT_RAM_11 = 256'h000036CCDCCC63000000F66667666F000000F66667666F000000F66666666F00;
defparam dpb_inst_1.INIT_RAM_12 = 256'h0000E66677666E0000007CCC0000010000003111111113000000CCCCCFCCCC00;
defparam dpb_inst_1.INIT_RAM_13 = 256'h00007CCCCCCCC7000000CCCCCDFFEC000000CCCCCDFFEC000000F66666666F00;
defparam dpb_inst_1.INIT_RAM_14 = 256'h00007CC0036CC7000000E66667666F0000007DDCCCCCC7000000F66667666F00;
defparam dpb_inst_1.INIT_RAM_15 = 256'h00006EFDDDCCCC000000136CCCCCCC0000007CCCCCCCCC000000311111157700;
defparam dpb_inst_1.INIT_RAM_16 = 256'h00003333333333000000FCC63108CF0000003111136666000000CC673376CC00;
defparam dpb_inst_1.INIT_RAM_17 = 256'h00F0000000000000000000000000C63100003000000003000000000137EC8000;
defparam dpb_inst_1.INIT_RAM_18 = 256'h00007CCCCC7000000000766666766E0000007CCC707000000000000000000133;
defparam dpb_inst_1.INIT_RAM_19 = 256'h07C07CCCCC7000000000F6666F66630000007CCCFC70000000007CCCC6300100;
defparam dpb_inst_1.INIT_RAM_1A = 256'h0000E66776666E00036600000000000000003111113011000000E66667666E00;
defparam dpb_inst_1.INIT_RAM_1B = 256'h00007CCCCC7000000000666666D000000000CDDDDFE000000000311111111300;
defparam dpb_inst_1.INIT_RAM_1C = 256'h00007C036C7000000000F66667D0000001007CCCCC7000000F66766666D00000;
defparam dpb_inst_1.INIT_RAM_1D = 256'h00006FDDDCC00000000013666660000000007CCCCCC000000000133333F33100;
defparam dpb_inst_1.INIT_RAM_1E = 256'h00000111171110000000FC631CF000000F007CCCCCC000000000C63336C00000;
defparam dpb_inst_1.INIT_RAM_1F = 256'h00000FCCC6310000000000000000D70000007111101117000000111110111100;
defparam dpb_inst_1.INIT_RAM_20 = 256'h00007CCC7070631000007CCCFC70310000007CCCCCC00C000070036CCCCC6300;
defparam dpb_inst_1.INIT_RAM_21 = 256'h000300366663000000007CCC7070363000007CCC7070136000007CCC70700C00;
defparam dpb_inst_1.INIT_RAM_22 = 256'h000031111130060000007CCCFC70136000007CCCFC700C0000007CCCFC706310;
defparam dpb_inst_1.INIT_RAM_23 = 256'h0000CCCFCC6303630000CCCFCC6310C000003111113013600000311111306310;
defparam dpb_inst_1.INIT_RAM_24 = 256'h00007CCCCC7063100000CCCCCFCC630000006DD737C000000000F666766F0631;
defparam dpb_inst_1.INIT_RAM_25 = 256'h00007CCCCCC0136000007CCCCCC0C73000007CCCCC70136000007CCCCC700C00;
defparam dpb_inst_1.INIT_RAM_26 = 256'h000011366666311000007CCCCCCCC0C000007CCCCCCC70C007007CCCCCC00C00;
defparam dpb_inst_1.INIT_RAM_27 = 256'h007D1111171111000000CCCCDCCFCCF000001117171366000000FE6666F66630;
defparam dpb_inst_1.INIT_RAM_28 = 256'h00007CCCCCC0631000007CCCCC706310000031111130310000007CCC70706310;
defparam dpb_inst_1.INIT_RAM_29 = 256'h000000000703663000000000070366300000CCCCDFFEC0D70000666666D0D700;
defparam dpb_inst_1.INIT_RAM_2A = 256'h003108D631CCCCC0000000000F00000000000CCCCF00000000007CCC63303300;
defparam dpb_inst_1.INIT_RAM_2B = 256'h000000D636D0000000000036D63000000000133311101100000039C631CCCCC0;
defparam dpb_inst_1.INIT_RAM_2C = 256'h11111111111111117D7D7D7D7D7D7D7DA5A5A5A5A5A5A5A54141414141414141;
defparam dpb_inst_1.INIT_RAM_2D = 256'h33333333F000000033333333F333333311111111F1F1111111111111F1111111;
defparam dpb_inst_1.INIT_RAM_2E = 256'h33333333F0F00000333333333333333333333333F0F3333311111111F1F00000;
defparam dpb_inst_1.INIT_RAM_2F = 256'h11111111F000000000000000F1F1111100000000F333333300000000F0F33333;
defparam dpb_inst_1.INIT_RAM_30 = 256'h111111111111111111111111F000000000000000F11111110000000011111111;
defparam dpb_inst_1.INIT_RAM_31 = 256'h3333333333333333111111111111111111111111F111111100000000F0000000;
defparam dpb_inst_1.INIT_RAM_32 = 256'h33333333F0F0000000000000F0F3333333333333333000000000000033333333;
defparam dpb_inst_1.INIT_RAM_33 = 256'h00000000F0F1111133333333F0F3333300000000F0F000003333333333333333;
defparam dpb_inst_1.INIT_RAM_34 = 256'h000000003333333333333333F000000011111111F0F0000000000000F3333333;
defparam dpb_inst_1.INIT_RAM_35 = 256'h33333333F3333333333333333000000011111111111000000000000011111111;
defparam dpb_inst_1.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFF111111111000000000000000F111111111111111F1F11111;
defparam dpb_inst_1.INIT_RAM_37 = 256'h000000000FFFFFFF0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFF0000000;
defparam dpb_inst_1.INIT_RAM_38 = 256'h00006666666F00000000CCCCCCCCCF000000CCCCCDCCC70000007DDDDD700000;
defparam dpb_inst_1.INIT_RAM_39 = 256'h0000111111D70000000C66766666000000007DDDDD7000000000FC63136CF000;
defparam dpb_inst_1.INIT_RAM_3A = 256'h00003666630131000000E6666CCC6300000036CCFCC630000000713666317000;
defparam dpb_inst_1.INIT_RAM_3B = 256'h0000CCCCCCCC700000001366676631000000C67FDD7000000000007DDD700000;
defparam dpb_inst_1.INIT_RAM_3C = 256'h000070013631000000007031000130000000F0011711000000000F00F00F0000;
defparam dpb_inst_1.INIT_RAM_3D = 256'h000000D70D700000000001107011000000007DDD111111111111111111111000;
defparam dpb_inst_1.INIT_RAM_3E = 256'h00001366E0000000000000010000000000000001100000000000000000036630;
defparam dpb_inst_1.INIT_RAM_3F = 256'h00000000000000000000077777770000000000000FC63D7000000000066666D0;

endmodule //Gowin_DPB_VGAFont
